module orgate(a,b,y);
input a,b;
output y;
or or1(y,a,b);
endmodule